/////////////////////////////////////////////
////     2Channel-Music-Synthesizer     /////
/////////////////////////////////////////////
/*****************************************************/
/*             KEY & SW List               			 */
/* BUTTON[1]: I2C reset                       		 */
/* BUTTON[2]: Demo Sound and Keyboard mode selection */
/* BUTTON[3]: Keyboard code Reset             		 */
/* BUTTON[4]: Keyboard system Reset                  */
/*****************************************************/

module synthesizer #(
parameter VOICES = 32,
parameter V_OSC = 4,				// number of oscilators pr. voice.
parameter O_ENVS = 2,				// number of envelope generators pr. oscilator.
parameter V_ENVS = V_OSC * O_ENVS,	// number of envelope generators  pr. voice.
parameter V_WIDTH = utils::clogb2(VOICES),
parameter O_WIDTH = utils::clogb2(V_OSC),
parameter OE_WIDTH = utils::clogb2(O_ENVS),
parameter E_WIDTH = O_WIDTH + OE_WIDTH,
AUD_BIT_DEPTH = 24
) (
// Clock
    input wire              data_clk,
    input wire              AUDIO_CLK,
// reset
    input wire              reset_n,
    input wire              trig,
// MIDI uart
    input wire              MIDI_Rx_DAT,
    output wire             midi_txd,

    input wire  [4:1]       button,
    output wire [VOICES-1:0] keys_on,
    output wire [VOICES-1:0] voice_free,

    output wire [AUD_BIT_DEPTH-1:0]  lsound_out,
    output wire [AUD_BIT_DEPTH-1:0]  rsound_out,

    output wire             xxxx_zero,

    input wire              io_reset_n,
    input wire              cpu_read,
    input wire              cpu_write,
    input wire              chipselect,
    input wire  [9:0]       address,
    output wire [31:0]      cpu_writedata,
    input wire  [31:0]      cpu_readdata,
    input wire              socmidi_read,
    input wire              socmidi_write,
    input wire              socmidi_cs,
    input wire  [2:0]       socmidi_addr,
    input wire  [7:0]       socmidi_data_in,
    output reg [7:0]        socmidi_data_out,
    output wire             run,
    input wire              uart_usb_sel
);

//-----		Registers		-----//
// io:

//    reg                 write_delay;
//    reg                 reg_w_act;
//    reg signed [7:0]    indata;
    wire [5:0]          cpu_sel;
    wire signed [7:0]   synth_data_out;
    wire signed [7:0]   synth_data_in;
//    wire w_act;
//    wire write_active;
    wire io_reset;
//    assign w_act = (cpu_write | write_delay);
//    assign write_active = (cpu_write | reg_w_act);
    assign io_reset = ~io_reset_n;

 //   assign synth_data_in = (!cpu_read && write_active) ? indata : 8'bz;
    assign synth_data_in = cpu_readdata[7:0];

addr_decoder #(.addr_width(3),.num_lines(6)) addr_decoder_inst
(
    .clk(data_clk) ,	// input  clk_sig
    .reset(io_reset) ,	// input  reset_sig
    .address(address[9:7]) ,	// input [addr_width-1:0] address_sig
    .sel(cpu_sel[5:0]) 	// output [num_lines:0] sel_sig
);

    wire data_DLY0, data_DLY1, data_DLY2, reg_DLY0, reg_DLY1, reg_DLY2;

    wire reg_reset_N;
    wire data_reset_N;
    wire reset_data_n;

    assign reg_reset_N = button[1] & reset_n;
    assign data_reset_N = button[2];

    wire reset_reg_N = reg_DLY2;
    assign reset_data_n = data_DLY1;

//---	Midi	---//
// inputs
    wire midi_rxd;
    assign midi_rxd = MIDI_Rx_DAT; // Direct to optocopler RS-232 port (fix it in in topfile)
//outputs
    wire midi_out_ready,midi_send_byte;
    wire [7:0] midi_out_data;
    wire byteready;
    wire [7:0] cur_status,midibyte_nr,midi_data_byte;

//---	Midi	Decoder ---//
    wire dataready;
    wire dec_sysex_data_patch_send;
// note events
    wire               	note_on;
    wire [V_WIDTH-1:0] 	cur_key_adr;
    wire [7:0]         	cur_key_val;
    wire [7:0]         	cur_vel_on;
    wire [7:0]         	cur_vel_off;
// from midi_controller_unit
    wire [13:0] 		pitch_val;
// from env gen

// inputs
// outputs
    wire octrl_cmd,prg_ch_cmd,pitch_cmd;
    wire[7:0] octrl,octrl_data,prg_ch_data;
    wire [V_WIDTH:0]	active_keys;
    wire 	off_note_error;

    wire ictrl_cmd;
    wire [7:0]ictrl, ictrl_data;

    wire HC_LCD_CLK, HC_VGA_CLOCK;

//    wire OSC_CLK;
    wire audio_pll_locked;

    wire [63:0] lvoice_out;
    wire [63:0] rvoice_out;

//---	Midi	Controllers unit ---//
    wire [6:0]	dec_addr;
    wire [6:0]	adr;
    wire [6:0]	dec_sel_bus;
    wire		env_sel	;
    wire		osc_sel;
    wire		m1_sel;
    wire		m2_sel;
    wire		com_sel;
    wire		read;
    wire		write;
    wire		sysex_data_patch_send;
    wire		dec_read_write;

    reg [3:0] midi_ch;
    reg [7:0] out_data;

addr_mux #(.addr_width(7),.num_lines(7)) addr_mux_inst
(
    .clk(data_clk) ,	// input  in_select_sig
    .dataready(dataready) ,	// input  in_select_sig
    .dec_syx(dec_sysex_data_patch_send) ,	// input  dec_syx_sig
    .cpu_and({chipselect,cpu_read}) ,	// input [1:0] cpu_and_sig
    .dec_addr(dec_addr) ,	// input [addr_width-1:0] dec_addr_sig
    .cpu_addr(address[6:0]) ,	// input [addr_width-1:0] cpu_addr_sig
    .cpu_sel({cpu_write,cpu_read,cpu_sel[5],cpu_sel[3:0]}) ,	// input [num_lines-1:0] cpu_sel_sig
    .dec_sel(dec_sel_bus) ,	// input [num_lines-1:0] dec_sel_sig
    .syx_out (sysex_data_patch_send),
    .addr_out(adr) ,	// output [addr_width-1:0] addr_out_sig
    .sel_out({write,read,com_sel,m2_sel,m1_sel,osc_sel,env_sel}) 	// output [num_lines-1:0] sel_out_sig
);


/** @brief write data
*/
    always@(negedge reg_reset_N or posedge data_clk)begin
        if(!reg_reset_N) begin
            midi_ch <= 4'h0;
        end else begin
            if(com_sel && write) begin
                if(adr == 2) midi_ch <= synth_data_in[3:0];
            end
        end
    end


/** @brief read data
*/
    always @(negedge data_clk) begin
        if(com_sel &&  read) begin
            if(adr == 2) out_data <= midi_ch;
        end
    end

    assign cpu_writedata = (com_sel && adr == 2) ? out_data : synth_data_out;

//    always @(posedge data_clk) begin
//        write_delay <= cpu_write;
//        reg_w_act <= w_act;
//    end
    
//    always @(posedge data_clk) begin
//        if (io_reset) begin
//            cpu_writedata[7:0] <= 8'b0;
//        end
//        else if (read) begin
//            cpu_writedata[7:0] <= (com_sel && adr == 2) ? out_data : synth_data_out;
//        end
//        else if    (write) begin
//            indata <= cpu_readdata[7:0];
//        end
//    end

////////////	Init Reset sig Gen	////////////
// system reset  //

reset_delay	reset_reg_delay_inst  (
    .iCLK(data_clk),
    .reset_reg_N(reg_reset_N),
    .oRST_0(reg_DLY0),
    .oRST_1(reg_DLY1),
    .oRST_2(reg_DLY2)
);

reset_delay	reset_data_delay_inst  (
    .iCLK(data_clk),
    .reset_reg_N(data_reset_N),
    .oRST_0(data_DLY0),
    .oRST_1(data_DLY1),
    .oRST_2(data_DLY2)
);

    // Sound clk gen //

synth_controller #(.VOICES(VOICES),.V_WIDTH(V_WIDTH)) synth_controller_inst(

    .reset_reg_N(reg_reset_N) ,
    .data_clk(data_clk) ,
    .socmidi_addr(socmidi_addr) ,
    .socmidi_data_in(socmidi_data_in) ,
    .socmidi_write(socmidi_write) ,
    .midi_rxd(midi_rxd) ,
    .midi_txd(midi_txd) ,
    .voice_free(voice_free) ,
    .midi_ch(midi_ch) ,

    .note_on(note_on) ,
    .keys_on(keys_on) ,
    .cur_key_adr(cur_key_adr) ,
    .cur_key_val(cur_key_val) ,
    .cur_vel_on(cur_vel_on) ,
    .cur_vel_off(cur_vel_off) ,
    .pitch_cmd(pitch_cmd) ,
    .octrl(octrl) ,
    .octrl_data(octrl_data) ,
    .prg_ch_cmd(prg_ch_cmd) ,
    .prg_ch_data(prg_ch_data) ,
// controller data bus
    .data_ready(dataready) ,
    .read_write (dec_read_write),
    .sysex_data_patch_send (dec_sysex_data_patch_send),
    .dec_addr(dec_addr) ,
    .synth_data_out (synth_data_out) ,
    .synth_data_in (synth_data_in) ,
    .dec_sel_bus( dec_sel_bus) ,
    .active_keys(active_keys) ,
    .uart_usb_sel(uart_usb_sel)
);


rt_controllers #(.VOICES(VOICES),.V_OSC(V_OSC)) rt_controllers_inst(
    .data_clk       ( data_clk ),
    .reset_data_N   ( reset_data_n ),
// from synth_controller
    .ictrl          ( octrl ),
    .ictrl_data     ( octrl_data ),
    .pitch_cmd      ( pitch_cmd ),
// outputs
    .pitch_val      ( pitch_val )
);

    //////////// Sound Generation /////////////

// 2CH Audio Sound output -- Audio Generater //
synth_engine #(.VOICES(VOICES),.V_OSC(V_OSC),.V_ENVS(V_ENVS),.V_WIDTH(V_WIDTH),.O_WIDTH(O_WIDTH),.OE_WIDTH(OE_WIDTH)) synth_engine_inst	(
// AUDIO CODEC //
    .AUDIO_CLK              ( AUDIO_CLK ),              // input
    .data_clk               ( data_clk ),
    .reset_reg_N            ( reg_reset_N ) ,           // input  reset_sig
    .reset_data_N           ( reg_reset_N ),
    .trig                   ( trig ),
    .lsound_out             ( lsound_out ),             //  Audio Raw Dat
    .rsound_out             ( rsound_out ),             //  Audio Raw Data
    .xxxx_zero              ( xxxx_zero) ,              // output  cycle complete signag
    // KEY //
    // -- Sound Control -- //
    //	to pitch control //
    .note_on                ( note_on ) ,               // input  note_on_sig
    .keys_on                ( keys_on ) ,               // input [VOICES-1:0] keys_on_sig
    .cur_key_adr            ( cur_key_adr ) ,           // input [V_WIDTH-1:0] cur_key_adr_sig
    .cur_key_val            ( cur_key_val ) ,           // input [7:0] cur_key_val_sig
    .cur_vel_on             ( cur_vel_on ) ,            // input [7:0] cur_vel_on_sig
    .cur_vel_off            ( cur_vel_off ) ,           // input [7:0] cur_vel_off_sig
// from midi_controller_unit
    .pitch_val              ( pitch_val ),
// controller data bus
    .write                  ( write) ,                  // input  write_sig
    .read                   ( read),                    // input read synth_data signal
    .sysex_data_patch_send  ( sysex_data_patch_send),   // input
    .adr                    ( adr) ,                    // input [6:0] adr_sig
    .synth_data_out         ( synth_data_out ) ,
    .synth_data_in          ( synth_data_in ) ,
    .env_sel                ( env_sel ) ,
    .osc_sel                ( osc_sel ) ,
    .m1_sel                 ( m1_sel ) ,
    .m2_sel                 ( m2_sel ) ,
    .com_sel                ( com_sel ),
// from env gen //
    .run                    ( run ),
    .voice_free             ( voice_free )              //output from envgen
);



endmodule
